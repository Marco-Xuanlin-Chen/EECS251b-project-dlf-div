module dummyDCO(
    input [7:0] row_sel_b,
    input [3:0] col_sel_b,
    output [2:0] stages
)

endmodule